module stimulus(clk, number);

input clk;
input [7:0] number;

endmodule
