module stimulus(clk, number);

input clk;
input [7:0] number [4:0];

endmodule
