module stimulus(clk, number[7:0]);
// module stimulus;

input clk;
input [7:0] number [4:0];

assign number[0] = 1'b1;

endmodule
