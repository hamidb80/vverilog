// module stimulus(clk, number[7:0]);
module stimulus;

// input clk;
input clk, load;
// input [7:0] number [4:0];
// assign number[0] = 1'b1;
// assign Word_Line_q1[1] = ~wrapout_s1[1] & phi1;

endmodule
