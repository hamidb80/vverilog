module stimulus(clk, number[7:0]);

input clk;
input [7:0] number [4:0];

endmodule
