module stimulus(clk, number[7:0]);

input clk;
input number;

endmodule
